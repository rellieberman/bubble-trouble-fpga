module startBitMap
(
        input	logic	clk,
        input	logic	resetN,
        input   logic	[10:0] offsetX,// offset from top left  position 
        input   logic	[10:0] offsetY,
        input	logic	InsideRectangle, //input that the pixel is within a bracket 

        output	logic	drawingRequest, //output that the pixel should be dispalyed 
        output	logic	[7:0] RGBout  //rgb value from the bitmap 
);

        localparam logic TRANSPARENT_ENCODING = 8'h00;// RGB value in the bitmap representing a transparent pixel 

        localparam  int OBJECT_WIDTH_X = 25;
        localparam  int OBJECT_HEIGHT_Y = 55;

        logic [0:OBJECT_HEIGHT_Y-1] [1*55-1:0] object_colors = {
        {55'b0000000000000000000000000000000000000000000000000000000},
        {55'b0000000000000000000000000000000000000000000000000000000},
        {55'b0000000000000000000000000000000000000000100000000000000},
        {55'b0000000000000000000000000000000000000000110000000000000},
        {55'b0000000000000000000000000000000000000000111000000000000},
        {55'b0000000011110011110011111001110001110000111110000000000},
        {55'b0000000011001011001011000011011011011000111111000000000},
        {55'b0000000010001010001011000011000011000000111111100000000},
        {55'b0000000011001011011011110001111001111000111111110000000},
        {55'b0000000011110011110011000000001100001100111111111000000},
        {55'b0000000010000010011011111001111001111000111111111100000},
        {55'b0000000000000000000000000000000000000000111111111111000},
        {55'b0000000000000000000000000000000000000000111111111111100},
        {55'b0000000000000000000000000000000000000000111111111111100},
        {55'b0000000000000000000000000000000000000000111111111111000},
        {55'b0001111001111110001110011111100011111100111111111110000},
        {55'b0011001000011000010010011000110000110000111111111100000},
        {55'b0011000000011000110011011000110000110000111111111000000},
        {55'b0001111000011000110011011001110000110000111111110000000},
        {55'b0000001100011000111111011111000000110000111111000000000},
        {55'b0010001100011000110011011011100000110000111110000000000},
        {55'b0011111100011000110011011001110000110000111100000000000},
        {55'b0000000000000000000000000000000000000000111000000000000},
        {55'b0000000000000000000000000000000000000000110000000000000},
        {55'b0000000000000000000000000000000000000000000000000000000}
        };
        
        always_ff@(posedge clk or negedge resetN)
        begin
            if(!resetN) begin
                RGBout <= 8'h00; 
            end
            else begin
                if (InsideRectangle && object_colors[offsetY>>1][offsetX>>1] )  // inside an external bracket 
                    RGBout <= 8'hFF; //black 
                else 
                    RGBout <= TRANSPARENT_ENCODING; // force color to transparent so it will not be displayed 
            end 
        end
        
    assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap  


endmodule

