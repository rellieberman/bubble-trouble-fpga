module charBitMap
    (
        input	logic	clk,
        input	logic	resetN,
        input   logic	[10:0] offsetX,// offset from top left  position 
        input   logic	[10:0] offsetY,
        input	logic	InsideRectangle, //input that the pixel is within a bracket 

        output	logic	drawingRequest, //output that the pixel should be dispalyed 
        output	logic	[7:0] RGBout  //rgb value from the bitmap 
    );
        
        localparam  int OBJECT_WIDTH_X = 32;
        localparam  int OBJECT_HEIGHT_Y = 20;

        localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 

        logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
        {8'h00, 8'h00, 8'h04, 8'h05, 8'h49, 8'h89, 8'hA9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hA9, 8'h89, 8'h65, 8'h44, 8'h00, 8'h04, 8'h05, 8'h05, },
        {8'h00, 8'h05, 8'h44, 8'hA9, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hED, 8'hED, 8'hC9, 8'hA9, 8'h44, 8'h05, 8'h00, },
        {8'h04, 8'h49, 8'hA4, 8'hA9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hA9, 8'hA4, 8'h45, 8'h00, },
        {8'h29, 8'hA9, 8'hC0, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC0, 8'hA9, 8'h25, },
        {8'h69, 8'hC9, 8'hC9, 8'hCD, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hA9, 8'hC9, 8'h49, },
        {8'h69, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hED, 8'h65, },
        {8'h49, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hED, 8'h45, },
        {8'h24, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'h24, },
        {8'h00, 8'hA9, 8'hE9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hE9, 8'h89, 8'h00, },
        {8'h00, 8'h49, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hA9, 8'hA9, 8'hA9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'h29, 8'h00, },
        {8'h00, 8'h04, 8'h49, 8'hC9, 8'hED, 8'hED, 8'h89, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h89, 8'hED, 8'hE9, 8'hC9, 8'h49, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h04, 8'h29, 8'hA9, 8'hC9, 8'h44, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h44, 8'hA9, 8'h89, 8'h24, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h04, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h09, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h29, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h29, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h04, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h00, 8'h05, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h04, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h05, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h04, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h04, 8'h00, 8'h00, 8'h00, },
        {8'h04, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h25, 8'h25, 8'h25, 8'h00, 8'h00, 8'h00, },
        {8'h00, 8'h00, 8'h25, 8'h24, 8'h25, 8'h24, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h25, 8'h24, 8'h24, 8'h68, 8'h48, 8'h09, 8'h00, 8'h00, },
        {8'h00, 8'h29, 8'h8C, 8'hB0, 8'h8C, 8'h68, 8'h68, 8'h68, 8'h68, 8'h29, 8'h29, 8'h68, 8'h68, 8'h68, 8'hAC, 8'hD0, 8'hD0, 8'hB0, 8'h29, 8'h00, },
        {8'h00, 8'h68, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h49, 8'h29, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h8C, 8'h04, }
        };

        // pipeline (ff) to get the pixel color from the array 	 

        always_ff@(posedge clk or negedge resetN)
        begin
            if(!resetN) begin
                RGBout <=	8'h00;
            end
            else begin
                if (InsideRectangle)  // inside an external bracket 
                    RGBout <= object_colors[offsetY][offsetX];	//get RGB from the colors table  
                else 
                    RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
            end 
        end

        // decide if to draw the pixel or not 
        assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap  

endmodule
